* C:\Users\mathias\Desktop\PED\LISTA_FINAL\lista_final.sch

* Schematics Version 9.1 - Web Update 1
* Mon Dec 10 17:41:55 2018



** Analysis setup **
.ac DEC 101 0.1 1e9
.OP 
.LIB "C:\Users\mathias\Desktop\PED\LISTA_FINAL\lista_final.lib"


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "lista_final.net"
.INC "lista_final.als"


.probe


.END
