* C:\Users\mathias\Desktop\PED\LISTA1\ex2\ex2.sch

* Schematics Version 9.1 - Web Update 1
* Fri Aug 03 16:29:05 2018



** Analysis setup **
.ac DEC 1000 0.1 1G


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "ex2.net"
.INC "ex2.als"


.probe


.END
