* C:\Users\mathias\Desktop\PED\LISTA2\ex2\ex2.sch

* Schematics Version 9.1 - Web Update 1
* Mon Aug 13 16:21:15 2018



** Analysis setup **
.tran 0ns 3m 0 1u
.LIB "C:\Users\mathias\Desktop\PED\LISTA2\ex2\ex2.lib"


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "ex2.net"
.INC "ex2.als"


.probe


.END
