* C:\Users\mathias\Desktop\PED\LISTA2\ex1\ex1.sch

* Schematics Version 9.1 - Web Update 1
* Mon Aug 13 18:20:30 2018



** Analysis setup **
.DC LIN V_V1 5 10 1 
.OP 
.LIB "C:\Users\mathias\Desktop\PED\LISTA2\ex1\ex1.lib"
.STMLIB "ex1.stl"


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "ex1.net"
.INC "ex1.als"


.probe


.END
