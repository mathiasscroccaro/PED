* C:\Users\mathias\Desktop\PED\LISTA1\sandbox2\Schematic1.sch

* Schematics Version 9.1 - Web Update 1
* Fri Sep 14 21:57:01 2018



** Analysis setup **
.ac DEC 101 0.1Hz 1GHz
.LIB "C:\Users\mathias\Desktop\PED\LISTA1\sandbox2\Schematic1.lib"


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic1.net"
.INC "Schematic1.als"


.probe


.END
