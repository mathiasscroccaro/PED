* C:\Users\mathias\Desktop\PED\LISTA1\ex2\ex2.sch

* Schematics Version 9.1 - Web Update 1
* Tue Oct 09 14:58:36 2018



** Analysis setup **
.ac DEC 1000 1 1G
.LIB "C:\Users\mathias\Desktop\PED\LISTA1\ex2\ex2.lib"


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "ex2.net"
.INC "ex2.als"


.probe


.END
