* C:\Users\mathias\Desktop\PED\LISTA1\ex3\ex3.sch

* Schematics Version 9.1 - Web Update 1
* Tue Oct 09 16:01:53 2018



** Analysis setup **
.ac DEC 100 0.1 1e9
.tran 0 10m 0 0.01m
.LIB "C:\Users\mathias\Desktop\PED\LISTA1\ex3\ex3.lib"


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "ex3.net"
.INC "ex3.als"


.probe


.END
