* C:\Users\mathias\Desktop\PED\LISTA1\ex1.sch

* Schematics Version 9.1 - Web Update 1
* Thu Jul 19 13:28:16 2018



** Analysis setup **
.DC LIN V_VGS 0 5 0.1 
.LIB "C:\Users\mathias\Desktop\PED\LISTA1\ex1.lib"


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "ex1.net"
.INC "ex1.als"


.probe


.END
